`timescale 1ns / 1ps
module inv_sbox(x,y,isbout);
input [0:3] x,y;
output reg [0:7] isbout;
always@(x,y)
begin
case({x,y})
8'h00:isbout =8'h52;
8'h01:isbout =8'h09;
8'h02:isbout =8'h6a;
8'h03:isbout =8'hd5;
8'h04:isbout =8'h30;
8'h05:isbout =8'h36;
8'h06:isbout =8'ha5;
8'h07:isbout =8'h38;
8'h08:isbout =8'hbf;
8'h09:isbout =8'h40;
8'h0a:isbout =8'ha3;
8'h0b:isbout =8'h9e;
8'h0c:isbout =8'h81;
8'h0d:isbout =8'hf3;
8'h0e:isbout =8'hd7;
8'h0f:isbout =8'hfb;
8'h10:isbout =8'h7c;
8'h11:isbout =8'he3;
8'h12:isbout =8'h39;
8'h13:isbout =8'h82;
8'h14:isbout =8'h9b;
8'h15:isbout =8'h2f;
8'h16:isbout =8'hff;
8'h17:isbout =8'h87;
8'h18:isbout =8'h34;
8'h19:isbout =8'h8e;
8'h1a:isbout =8'h43;
8'h1b:isbout =8'h44;
8'h1c:isbout =8'hc4;
8'h1d:isbout =8'hde;
8'h1e:isbout =8'he9;
8'h1f:isbout =8'hcb;
8'h20:isbout =8'h54;
8'h21:isbout =8'h7b;
8'h22:isbout =8'h94;
8'h23:isbout =8'h32;
8'h24:isbout =8'ha6;
8'h25:isbout =8'hc2;
8'h26:isbout =8'h23;
8'h27:isbout =8'h3d;
8'h28:isbout =8'hee;
8'h29:isbout =8'h4c;
8'h2a:isbout =8'h95;
8'h2b:isbout =8'h0b;
8'h2c:isbout =8'h42;
8'h2d:isbout =8'hfa;
8'h2e:isbout =8'hc3;
8'h2f:isbout =8'h4e;
8'h30:isbout =8'h08;
8'h31:isbout =8'h2e;
8'h32:isbout =8'ha1;
8'h33:isbout =8'h66;
8'h34:isbout =8'h28;
8'h35:isbout =8'hd9;
8'h36:isbout =8'h24;
8'h37:isbout =8'hb2;
8'h38:isbout =8'h76;
8'h39:isbout =8'h5b;
8'h3a:isbout =8'ha2;
8'h3b:isbout =8'h49;
8'h3c:isbout =8'h6d;
8'h3d:isbout =8'h8b;
8'h3e:isbout =8'hd1;
8'h3f:isbout =8'h25;
8'h40:isbout =8'h72;
8'h41:isbout =8'hf8;
8'h42:isbout =8'hf6;
8'h43:isbout =8'h64;
8'h44:isbout =8'h86;
8'h45:isbout =8'h68;
8'h46:isbout =8'h98;
8'h47:isbout =8'h16;
8'h48:isbout =8'hd4;
8'h49:isbout =8'ha4;
8'h4a:isbout =8'h5c;
8'h4b:isbout =8'hcc;
8'h4c:isbout =8'h5d;
8'h4d:isbout =8'h65;
8'h4e:isbout =8'hb6;
8'h4f:isbout =8'h92;
8'h50:isbout =8'h6c;
8'h51:isbout =8'h70;
8'h52:isbout =8'h48;
8'h53:isbout =8'h50;
8'h54:isbout =8'hfd;
8'h55:isbout =8'hed;
8'h56:isbout =8'hb9;
8'h57:isbout =8'hda;
8'h58:isbout =8'h5e;
8'h59:isbout =8'h15;
8'h5a:isbout =8'h46;
8'h5b:isbout =8'h57;
8'h5c:isbout =8'ha7;
8'h5d:isbout =8'h8d;
8'h5e:isbout =8'h9d;
8'h5f:isbout =8'h84;
8'h60:isbout =8'h90;
8'h61:isbout =8'hd8;
8'h62:isbout =8'hab;
8'h63:isbout =8'h00;
8'h64:isbout =8'h8c;
8'h65:isbout =8'hbc;
8'h66:isbout =8'hd3;
8'h67:isbout =8'h0a;
8'h68:isbout =8'hf7;
8'h69:isbout =8'he4;
8'h6a:isbout =8'h58;
8'h6b:isbout =8'h05;
8'h6c:isbout =8'hb8;
8'h6d:isbout =8'hb3;
8'h6e:isbout =8'h45;
8'h6f:isbout =8'h06;
8'h70:isbout =8'hd0;
8'h71:isbout =8'h2c;
8'h72:isbout =8'h1e;
8'h73:isbout =8'h8f;
8'h74:isbout =8'hca;
8'h75:isbout =8'h3f;
8'h76:isbout =8'h0f;
8'h77:isbout =8'h02;
8'h78:isbout =8'hc1;
8'h79:isbout =8'haf;
8'h7a:isbout =8'hbd;
8'h7b:isbout =8'h03;
8'h7c:isbout =8'h01;
8'h7d:isbout =8'h13;
8'h7e:isbout =8'h8a;
8'h7f:isbout =8'h6b;
8'h80:isbout =8'h3a;
8'h81:isbout =8'h91;
8'h82:isbout =8'h11;
8'h83:isbout =8'h41;
8'h84:isbout =8'h4f;
8'h85:isbout =8'h67;
8'h86:isbout =8'hdc;
8'h87:isbout =8'hea;
8'h88:isbout =8'h97;
8'h89:isbout =8'hf2;
8'h8a:isbout =8'hcf;
8'h8b:isbout =8'hce;
8'h8c:isbout =8'hf0;
8'h8d:isbout =8'hb4;
8'h8e:isbout =8'he6;
8'h8f:isbout =8'h73;
8'h90:isbout =8'h96;
8'h91:isbout =8'hac;
8'h92:isbout =8'h74;
8'h93:isbout =8'h22;
8'h94:isbout =8'he7;
8'h95:isbout =8'had;
8'h96:isbout =8'h35;
8'h97:isbout =8'h85;
8'h98:isbout =8'he2;
8'h99:isbout =8'hf9;
8'h9a:isbout =8'h37;
8'h9b:isbout =8'he8;
8'h9c:isbout =8'h1c;
8'h9d:isbout =8'h75;
8'h9e:isbout =8'hdf;
8'h9f:isbout =8'h6e;
8'ha0:isbout =8'h47;
8'ha1:isbout =8'hf1;
8'ha2:isbout =8'h1a;
8'ha3:isbout =8'h71;
8'ha4:isbout =8'h1d;
8'ha5:isbout =8'h29;
8'ha6:isbout =8'hc5;
8'ha7:isbout =8'h89;
8'ha8:isbout =8'h6f;
8'ha9:isbout =8'hb7;
8'haa:isbout =8'h62;
8'hab:isbout =8'h0e;
8'hac:isbout =8'haa;
8'had:isbout =8'h18;
8'hae:isbout =8'hbe;
8'haf:isbout =8'h1b;
8'hb0:isbout =8'hfc;
8'hb1:isbout =8'h56;
8'hb2:isbout =8'h3e;
8'hb3:isbout =8'h4b;
8'hb4:isbout =8'hc6;
8'hb5:isbout =8'hd2;
8'hb6:isbout =8'h79;
8'hb7:isbout =8'h20;
8'hb8:isbout =8'h9a;
8'hb9:isbout =8'hdb;
8'hba:isbout =8'hc0;
8'hbb:isbout =8'hfe;
8'hbc:isbout =8'h78;
8'hbd:isbout =8'hcd;
8'hbe:isbout =8'h5a;
8'hbf:isbout =8'hf4;
8'hc0:isbout =8'h1f;
8'hc1:isbout =8'hdd;
8'hc2:isbout =8'ha8;
8'hc3:isbout =8'h33;
8'hc4:isbout =8'h88;
8'hc5:isbout =8'h07;
8'hc6:isbout =8'hc7;
8'hc7:isbout =8'h31;
8'hc8:isbout =8'hb1;
8'hc9:isbout =8'h12;
8'hca:isbout =8'h10;
8'hcb:isbout =8'h59;
8'hcc:isbout =8'h27;
8'hcd:isbout =8'h80;
8'hce:isbout =8'hec;
8'hcf:isbout =8'h5f;
8'hd0:isbout =8'h60;
8'hd1:isbout =8'h51;
8'hd2:isbout =8'h7f;
8'hd3:isbout =8'ha9;
8'hd4:isbout =8'h19;
8'hd5:isbout =8'hb5;
8'hd6:isbout =8'h4a;
8'hd7:isbout =8'h0d;
8'hd8:isbout =8'h2d;
8'hd9:isbout =8'he5;
8'hda:isbout =8'h7a;
8'hdb:isbout =8'h9f;
8'hdc:isbout =8'h93;
8'hdd:isbout =8'hc9;
8'hde:isbout =8'h9c;
8'hdf:isbout =8'hef;
8'he0:isbout =8'ha0;
8'he1:isbout =8'he0;
8'he2:isbout =8'h3b;
8'he3:isbout =8'h4d;
8'he4:isbout =8'hae;
8'he5:isbout =8'h2a;
8'he6:isbout =8'hf5;
8'he7:isbout =8'hb0;
8'he8:isbout =8'hc8;
8'he9:isbout =8'heb;
8'hea:isbout =8'hbb;
8'heb:isbout =8'h3c;
8'hec:isbout =8'h83;
8'hed:isbout =8'h53;
8'hee:isbout =8'h99;
8'hef:isbout =8'h61;
8'hf0:isbout =8'h17;
8'hf1:isbout =8'h2b;
8'hf2:isbout =8'h04;
8'hf3:isbout =8'h7e;
8'hf4:isbout =8'hba;
8'hf5:isbout =8'h77;
8'hf6:isbout =8'hd6;
8'hf7:isbout =8'h26;
8'hf8:isbout =8'he1;
8'hf9:isbout =8'h69;
8'hfa:isbout =8'h14;
8'hfb:isbout =8'h63;
8'hfc:isbout =8'h55;
8'hfd:isbout =8'h21;
8'hfe:isbout =8'h0c;
8'hff:isbout =8'h7d;
endcase
end
endmodule
